module rom(address,data);
input [8:0] address; //needs to be changed
output [38:0] data;	//needs to be changed
reg [38:0] array[511:0];	//needs to be changed
always @*
begin
//array[] = 39'b000000000_000_00010100_0000000000_00000_0000;

//nop
array[0]= 39'b000000001_000_00000000_0000000000_00000_0000;

//fetch and decode
array[1] = 39'b000000010_000_00000000_0000000000_00001_0000;
array[2] = 39'b000000011_000_00000000_0000001000_00000_0000;
array[3] = 39'b000000000_100_00110101_0000000100_00000_0110;

//bipush
array[16] = 39'b000010001_000_00110101_0000100001_00001_0011;
array[17] = 39'b000010010_000_00010100_0000001000_00000_0000;
array[18] = 39'b100010001_000_00010100_0000010010_00000_0101;
array[273] = 39'b100010010_000_00110101_0000000100_00100_0110;
array[274] = 39'b000000001_000_00010100_0000000000_01000_0000;

//ldc_w
array[19] = 39'b000010100_000_00110101_0000000100_00001_0110;
array[20] = 39'b100010011_000_00010100_0000001000_00000_0000;
array[275] = 39'b100010100_000_01010100_1000000000_00001_1101;
array[276] = 39'b100011111_000_00010100_0000001000_00000_0000;
array[287] = 39'b100100000_000_00011100_1000000000_00000_0101;
array[288] = 39'b100100001_000_00111100_0000000001_00000_0001;
array[289] = 39'b100100010_000_00110101_0000100001_00010_0011;
array[290] = 39'b100100011_000_00010100_0000000010_10000_0000;
array[291] = 39'b100100100_000_00110101_0000000100_00100_0110;
array[292] = 39'b000000001_000_00010100_0000010000_01000_0111;

//iload
array[21] = 39'b000010110_000_00010100_1000000000_00001_0010;
array[22] = 39'b000010111_000_00010100_0000001000_00000_0000;
array[23] = 39'b000011000_000_00111100_0000000001_00000_1101;
array[24] = 39'b000011001_000_00110101_0000100001_00010_0011;
array[25] = 39'b000011010_000_00010100_0000000010_10000_0000;
array[26] = 39'b000011011_000_00110101_0000000100_00100_0110;
array[27] = 39'b000000001_000_00010100_0000010000_01000_0111;

//istore
array[54] = 39'b000110111_000_00010100_1000000000_00001_0010;
array[55] = 39'b000111000_000_00010100_0000001000_00000_0000;
array[56] = 39'b000111001_000_00010100_0000000010_00000_0100;
array[57] = 39'b000111010_000_00111100_0000000001_00000_1101;
array[58] = 39'b000111011_000_00110110_0000100001_00100_0011;
array[59] = 39'b000111100_000_00010100_0000000000_01000_0000;
array[60] = 39'b000111101_000_00110101_0000000100_00010_0110;
array[61] = 39'b000111110_000_00010100_0000000000_10000_0000;
array[62] = 39'b000000001_000_00010100_0000010000_00000_0111;

//pop
array[87] = 39'b001011000_000_00110110_0000100001_00000_0011;
array[88] = 39'b000000000_000_00010100_0000000000_00010_0000;
array[271] = 39'b100001111_000_00010100_0000000010_00000_0000;
array[272] = 39'b000000001_000_00010100_0000010000_00000_0111;

//dup
array[89] = 39'b001011010_000_00110101_0000100001_00000_0011;
array[90] = 39'b001011011_000_00010100_0000000010_00000_0000;
array[91] = 39'b001011100_000_00010100_0000000000_00100_0000;
array[92] = 39'b000000001_000_00010100_0000000000_01000_0000;

//swap
array[95] = 39'b100001001_000_00110110_0000000001_00010_0011;
array[265] = 39'b100001010_000_00010100_0000000011_10000_0011;
array[266] = 39'b100001011_000_00010100_0100000000_00100_0111;
array[267] = 39'b100001100_000_00010100_0000000010_01000_0100;
array[268] = 39'b100001101_000_00110110_0000000001_00000_0011;
array[269] = 39'b100001110_000_00010100_0000010000_00100_0000;
array[270] = 39'b000000001_000_00010100_0000000000_01000_0000;

//iadd
array[96] = 39'b001100001_000_00110110_0000100001_00000_0011;
array[97] = 39'b001100010_000_00010100_1000000000_00010_0100;
array[98] = 39'b001100011_000_00010100_0000000010_10000_0000;
array[99] = 39'b100000000_000_00111100_0000010010_00000_0111;
array[256] = 39'b100000001_000_00010100_0000000000_00100_0000;
array[257] = 39'b000000001_000_00010100_0000000000_01000_0000;

//isub
array[100] = 39'b001100101_000_00110110_0000100001_00000_0011;
array[101] = 39'b001100110_000_00010100_1000000000_00010_0100;
array[102] = 39'b001100111_000_00010100_0000000010_10000_0000;
array[103] = 39'b001101000_000_00111111_0000010010_00000_0111;
array[104] = 39'b001101001_000_00010100_0000000000_00100_0000;
array[105] = 39'b000000001_000_00010100_0000000000_01000_0000;

//iand
array[126] = 39'b001111111_000_00110110_0000100001_00000_0011;
array[127] = 39'b100000010_000_00010100_1000000000_00010_0100;
array[258] = 39'b100000011_000_00010100_0000000010_10000_0000;
array[259] = 39'b100000100_000_00001100_0000010010_00000_0111;
array[260] = 39'b100000101_000_00010100_0000000000_00100_0000;
array[261] = 39'b000000001_000_00010100_0000000000_01000_0000;

//ior
array[128] = 39'b010000001_000_00110110_0000100001_00000_0011;
array[129] = 39'b010000010_000_00010100_1000000000_00010_0100;
array[130] = 39'b010000011_000_00010100_0000000010_10000_0000;
array[131] = 39'b100000110_000_00011100_0000010010_00000_0111;
array[262] = 39'b100000111_000_00010100_0000000000_00100_0000;
array[263] = 39'b000000001_000_00010100_0000000000_01000_0000;

//iinc
array[132] = 39'b010000101_000_00110101_0000000100_00001_0110;
array[133] = 39'b010000110_000_00010100_1000001000_00000_0010;
array[134] = 39'b010000111_000_00111100_0000000001_00001_1101;
array[135] = 39'b010001000_000_00010100_0000001000_00010_0000;
array[136] = 39'b010001001_000_00010100_0000000010_10000_0000;
array[137] = 39'b010001010_000_00010100_1000000000_00000_0111;
array[138] = 39'b010001011_000_00111100_0000000010_00000_0101;
array[139] = 39'b010001100_000_00110101_0000000100_00100_0110;
array[140] = 39'b000000001_000_00010100_0000000000_01000_0000;

//ifeq
array[153] = 39'b010011010_000_00110110_0000100001_00000_0011;
array[154] = 39'b100011011_000_00010100_0100000000_00010_0100;
array[283] = 39'b100011100_000_00010100_0000000010_10000_0000;
array[284] = 39'b100011101_000_00010100_0000010000_00000_0111;
array[285] = 39'b011111010_001_10010100_0000000000_00000_0000;

//iflt
array[155] = 39'b010011100_000_00110110_0000100001_00000_0011;
array[156] = 39'b010011101_000_00010100_0100000000_00010_0100;
array[157] = 39'b010011110_000_00010100_0000000010_10000_0000;
array[158] = 39'b100011110_000_00010100_0000010000_00000_0111;
array[286] = 39'b011111010_010_10010100_0000000000_00000_0000;

//if_icmpeq
array[159] = 39'b010100000_000_00110110_0000100001_00000_0011;
array[160] = 39'b010100001_000_00110110_0000100001_00010_0011;
array[161] = 39'b010100010_000_00010100_0100000010_10000_0100;
array[162] = 39'b010100011_000_00010100_1000000000_00010_0111;
array[163] = 39'b010100100_000_00010100_0000000010_10000_0000;
array[164] = 39'b010100101_000_00010100_0000010000_00000_0111;
array[165] = 39'b011111010_001_10111111_0000000000_00000_0000;

//True
array[506] = 39'b010101000_000_00110110_0100000000_00000_0110;

//False
array[250] = 39'b011111011_000_00110101_0000000100_00000_0110;
array[251] = 39'b000000001_000_00110101_0000000100_00000_0110;


//goto
array[167] = 39'b010101000_000_00110110_0100000000_00000_0110;
array[168] = 39'b010101001_000_00110101_0000000100_00001_0110;
array[169] = 39'b010101010_000_01010100_1000000000_00001_0101;
array[170] = 39'b010101011_000_00010100_0000001000_00000_0000;
array[171] = 39'b100001000_000_00011100_1000000000_00000_1101;
array[264] = 39'b000000001_000_00111100_0000000100_00000_0000;

//ireturn
array[172] = 39'b010101101_000_00010100_0000100001_00000_0010;
array[173] = 39'b010101110_000_00010100_0000000000_00010_0000;
array[174] = 39'b010101111_000_00010100_0000000010_10000_0000;
array[175] = 39'b010110000_000_00010100_0001000001_00000_0111;
array[176] = 39'b010110001_000_00010100_0000000000_00010_0000;
array[177] = 39'b010110010_000_00010100_0000000010_10000_0000;
array[178] = 39'b010110011_000_00110101_0000000001_00000_0010;
array[179] = 39'b010110100_000_00010100_0000000100_00010_0111;
array[180] = 39'b010110101_000_00010100_0000000011_10000_0011;
array[181] = 39'b100100101_000_00010100_0001000000_00000_0111;
array[293] = 39'b100100110_000_00010100_0000000010_00000_0100;
array[294] = 39'b100100111_000_00010100_0000000000_00100_0000;
array[295] = 39'b000000001_000_00010100_0000000000_01000_0000;

//invokevirtual
array[182] = 39'b010110111_000_00110101_0000000100_00001_0110;
array[183] = 39'b010111000_000_00010100_0000001000_00000_0000;
array[184] = 39'b010111001_000_01010100_1000000000_00001_0101;
array[185] = 39'b010111010_000_00010100_0000001000_00000_0000;
array[186] = 39'b010111011_000_00011100_1000000000_00000_1101;
array[187] = 39'b010111100_000_00111100_0000000001_00000_0001;
array[188] = 39'b010111101_000_00110101_0100000000_00010_0110;
array[189] = 39'b010111110_000_00010100_0000000010_10000_0000;
array[190] = 39'b010111111_000_00010100_0000000100_00000_0111;
array[191] = 39'b011000000_000_00110101_0000000100_00001_0110;
array[192] = 39'b011000001_000_00010100_0000001000_00000_0000;
array[193] = 39'b011000010_000_01010100_1000000000_00001_0101;
array[194] = 39'b011000011_000_00010100_0000001000_00000_0000;
array[195] = 39'b100101000_000_00110101_0000000100_00000_0110;
array[296] = 39'b100101001_000_00011100_1000000000_00001_1101;
array[297] = 39'b100101010_000_00010100_0000001000_00000_0000;
array[298] = 39'b100101011_000_00111111_0000010000_00000_0011;
array[299] = 39'b100101100_000_00110101_0000010001_00000_0100;
array[300] = 39'b100101101_000_00110101_0000000100_00001_0110;
array[301] = 39'b100101110_000_00010100_0000001000_00000_0000;
array[302] = 39'b100101111_000_01010100_1000000000_00001_0101;
array[303] = 39'b100110000_000_00010100_0000001000_00000_0000;
array[304] = 39'b100110001_000_00011100_1000000000_00000_1101;
array[305] = 39'b100110010_000_00111101_0000000010_00000_0011;
array[306] = 39'b100110011_000_00010100_0000100001_00100_0111;
array[307] = 39'b100110100_000_00010100_0000000000_01000_0000;
array[308] = 39'b100110101_000_00010100_0000000010_00000_0000;
array[309] = 39'b100111100_000_00110101_0000000100_00100_0110;
array[316] = 39'b100111101_000_00010100_0000000000_01000_0000;
array[317] = 39'b100111110_000_00110101_0000100001_00000_0011;
array[318] = 39'b100111111_000_00010100_0000000010_00001_0010;
array[319] = 39'b101000000_000_00010100_0000001000_00100_0000;
array[320] = 39'b000000001_000_00010100_0001000000_01000_0100;

//wide
array[196] = 39'b011000101_000_00110101_0000000100_00001_0110;
array[197] = 39'b011000110_000_00010100_0000001000_00000_0000;
array[198] = 39'b100000000_100_00010100_0000000000_00000_0000;

//wide_iload
array[277] = 39'b100010110_000_00110101_0000000100_00001_0110;
array[278] = 39'b100010111_000_00010100_0000001000_00000_0000;
array[279] = 39'b100011000_000_01010100_1000000000_00001_0101;
array[280] = 39'b100011001_000_00010100_0000001000_00000_0000;
array[281] = 39'b100011010_000_00011100_1000000000_00000_1101;
array[282] = 39'b000011000_000_00111100_0000000001_00000_0010;

//wide_istore
array[310] = 39'b100110111_000_00110101_0000000100_00001_0110;
array[311] = 39'b100111000_000_00010100_0000001000_00000_0000;
array[312] = 39'b100111001_000_01010100_1000000000_00001_0101;
array[313] = 39'b100111010_000_00010100_0000001000_00000_0000;
array[314] = 39'b100111011_000_00011100_1000000000_00000_1101;
array[315] = 39'b000111010_000_00111100_0000000001_00000_0010;

//wide_iinc
array[388] = 39'b110000101_000_00110101_0000000100_00001_0110;
array[389] = 39'b110000110_000_00010100_0000001000_00000_0000;
array[370] = 39'b110000111_000_01010100_1000000000_00000_0101;
array[371] = 39'b110001000_000_00110101_0000000100_00001_0110;
array[372] = 39'b110001001_000_00010100_0000001000_00000_0000;
array[373] = 39'b110001010_000_00011100_1000000000_00000_1101;
array[374] = 39'b010001000_000_00111100_0000000001_00000_0010;

end
assign data=array[address];
endmodule
